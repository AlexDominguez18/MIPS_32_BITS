
module MIPS_32_BITS(
	input A,
	output B
);

endmodule 